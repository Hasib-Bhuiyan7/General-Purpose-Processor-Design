library verilog;
use verilog.vl_types.all;
entity Processor_vlg_vec_tst is
end Processor_vlg_vec_tst;
