LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY for4To16decoder IS
	PORT (w  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0) ;
			En : IN  STD_LOGIC ;
			Y:  OUT STD_LOGIC_VECTOR(0 TO 15))  ;
		
END for4To16decoder ;

ARCHITECTURE Behavior OF for4To16decoder IS
	SIGNAL Enw : STD_LOGIC_VECTOR(4 DOWNTO 0) ;
BEGIN
	Enw <= En & w(3)&w(2)&w(1)&w(0);
	WITH Enw SELECT --[Enw + y] => ["Enw"+"0000"]
	Y <=    
	  "0000000000000001" WHEN "10000",
	  "0000000000000010" WHEN "10001",
	  "0000000000000100" WHEN "10010",
	  "0000000000001000" WHEN "10011",
	  "0000000000010000" WHEN "10100",
	  "0000000000100000" WHEN "10101",
	  "0000000001000000" WHEN "10110",
	  "0000000010000000" WHEN "10111",
	  "0000000100000000" WHEN "11000",
	  "0000000000000001" WHEN OTHERS;
			
		
END Behavior ;